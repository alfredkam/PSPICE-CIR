** PSPICE = power supply design (fig2) **

** +vdd +55v @ V(6,0) , -vdd -55v @(16,0)

* 1 mA Diode Model 
*
.model 1mA_diode D   (Is=100pA n=1.679 )

* 1N5402 2A Rectifier Diode <data sheet> (used as zener to regulate the voltage)
*
.model D1N5402 D (
+ Is=11.5f Rs=8.254m Ikf=3.87 N=1 Xti=3 Eg=1.11 Cjo=130.4p
+ M=.3758 Vj=.75 Fc=.5 Isr=61.19u Nr=2 )

.subckt zener_diode 1 2
* connections: | |
* anode |
* cathode
Dforward 1 2 1mA_diode
Dreverse 2 4 1mA_diode
Vz0 4 3 DC 4.9V 
Rz 1 3 10
* diode model statements
.model 1mA_diode D (Is=100pA n=1.679 )
.model ideal_diode D (Is=100pA n=0.01 )
.ends zener_diode

** main circuit **
* ac line voltage 
* positive vdd

Vac1 9 0 sin (0 120V 60Hz 0 0)
Rg1 9 1 100

* transformer section center tap
Lp1 1 0 4.57
Ls1 2 0 1
Kxfrmr1 Lp1 Ls1 0.99999


D1 2 6 1mA_diode
C1 0 6 500uF
Rs1 6 7 225k
XZ1 7 0 zener_diode

* negative vdd
Vac2 10 0 sin (0 120V 60Hz 0 0)
Rg2 10 11 100

* transformer section center tap
Lp2 11 0 4.57
Ls2 12 0 1
Kxfrmr2 Lp2 Ls2 0.99999


D2 16 12 1mA_diode
C2 0 16 500uF
Rs2 16 17 225k
XZ2 17 0 zener_diode




** analysis requests
.OPTIONS ITL5=0
.TRAN 0.5ms 5s 0ms 0.5ms UIC

** output requests
.PROBE
.END
 
