** PSPICE = power supply design (fig2) **

** PS +VDD +55V @ V(6,0), -VDD -55V @ V(16,0) 
** right speaker 10Vpp ~ AC 5V @ V(23,0)
** left speaker 10Vpp ~ AC 5V @ V(25,0)

** models
* 1 mA Diode Model 
*
.model 1mA_diode D   (Is=100pA n=1.679 )

* 1N5402 2A Rectifier Diode <data sheet> (used as zener to regulate the voltage)
*
.model D1N5402 D (
+ Is=11.5f Rs=8.254m Ikf=3.87 N=1 Xti=3 Eg=1.11 Cjo=130.4p
+ M=.3758 Vj=.75 Fc=.5 Isr=61.19u Nr=2 )

.subckt zener_diode 1 2
* connections: | |
* anode |
* cathode
Dforward 1 2 1mA_diode
Dreverse 2 4 1mA_diode
Vz0 4 3 DC 4.9V 
Rz 1 3 10
* diode model statements
.model 1mA_diode D (Is=100pA n=1.679 )
.model ideal_diode D (Is=100pA n=0.01 )
.ends zener_diode

* 741 Op Amp Model <data sheet>
*
* UA741 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 07/05/89 AT 09:09
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT UA741    1 2 3 4 5
*
  C1   11 12 4.664E-12
  C2    6  7 20.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 10.61E6 -10E6 10E6 10E6 -10E6
  GA 6  0 11 12 137.7E-6
  GCM 0  6 10 99 2.574E-9
  IEE  10  4 DC 10.16E-6
  HLIM 90  0 VLIM 1K
  Q1   11  2 13 QX
  Q2   12  1 14 QX
  R2    6  9 100.0E3
  RC1   3 11 7.957E3
  RC2   3 12 7.957E3
  RE1  13 10 2.740E3
  RE2  14 10 2.740E3
  REE  10 99 19.69E6
  RO1   8  5 150
  RO2   7 99 150
  RP    3  4 18.11E3
  VB    9  0 DC 0
  VC 3 53 DC 2.600
  VE   54  4 DC 2.600
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL QX NPN(IS=800.0E-18 BF=62.50)
.ENDS

** main circuit **
* ac line voltage 
* positive vdd

Vac1 9 0 AC 1 sin(0 120V 60Hz 0 0)
Rg1 9 1 100

* transformer section center tap
Lp1 1 0 4.57
Ls1 2 0 1
Kxfrmr1 Lp1 Ls1 0.99999


D1 2 6 1mA_diode
C1 0 6 500uF
Rs1 6 7 225k
XZ1 7 0 zener_diode

* negative vdd
Vac2 10 0 AC 1 sin(0 120V 60Hz 0 0)
Rg2 10 11 100

* transformer section center tap
Lp2 11 0 4.57
Ls2 12 0 1
Kxfrmr2 Lp2 Ls2 0.99999


D2 16 12 1mA_diode
C2 0 16 500uF
Rs2 16 17 225k
XZ2 17 0 zener_diode

*********** ipod ****

Vac 21 0 AC 1 sin(0 250mv 60Hz 0 0)
Ripod 21 22 100

Xop1 22 24 6 16 23 UA741
R11 0 24 100
R12 24 23 2K
Rspeaker1 23 0 100K

Xop2 22 26 6 16 25 UA741
R21 0 26 100
R22 26 25 2K
Rspeaker2 25 0 100K



** analysis requests
.OPTIONS ITL5=0
.TRAN 0.5ms 5s 0ms 0.5ms UIC

** output requests
.PROBE
.END
 
